module viscord

// todo: http discord api calls